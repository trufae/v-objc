module uikit
