module objc

fn C.ivar_getName(Id) Id
fn C.ivar_getTypeEncoding(Id) Id
fn C.ivar_getOffset(Id) Id
