module objc

/*
    "protocol_getName": ['pointer', ['pointer']],
    "protocol_copyMethodDescriptionList": ['pointer', ['pointer', 'bool', 'bool', 'pointer']],
    "protocol_copyPropertyList": ['pointer', ['pointer', 'pointer']],
    "protocol_copyProtocolList": ['pointer', ['pointer', 'pointer']],
    "protocol_addProtocol": ['void', ['pointer', 'pointer']],
    "protocol_addMethodDescription": ['void', ['pointer', 'pointer', 'pointer', 'bool', 'bool']],
*/
