module objc
/*
    "property_getName": ['pointer', ['pointer']],
    "property_copyAttributeList": ['pointer', ['pointer', 'pointer']],
*/
